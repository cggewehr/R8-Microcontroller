--------------------------------------------------------------------------------
-- Project     : R8Gen
--------------------------------------------------------------------------------
-- File        : R8_PKG.vhd
-- Authors     : Carlos Gewehr(carlos.gewehr@ecomp.ufsm.br), 
--               Emilio Ferreira(emilio.ferreira@ecomp.ufsm.br)
-- Standard    : VHDL-1993
--------------------------------------------------------------------------------
-- Description : Template for software generated R8_pkg file, which contains 
--              configuration values for the R8 processor.
--------------------------------------------------------------------------------
-- Changelog   : v0.01 - Gewehr: Initial commit, defines project template
--------------------------------------------------------------------------------


package R8_PKG is

	-- R8 processor instructions. To be autogenerated by software
	type R8Instruction_t is (

		-- Basic Instructions
		ADD, SUB, AAND, OOR, XXOR, ADDI, SUBI, NNOT,
        SL0, SL1, SR0, SR1,
        LDL, LDH, LD, ST, LDSP, POP, PUSH,
        JMPR, JMPNR, JMPZR, JMPCR, JMPVR,  -- JUMP_R
        JMP, JMPN, JMPZ, JMPC, JMPV,       -- JUMP_A
        JMPD, JMPND, JMPZD, JMPCD, JMPVD,  -- JUMP_D
        JSRR, JSR, JSRD,
        NOP, HALT, RTS, INVALID

        -- Multiplication and Division
        MUL, DIV, MFH, MFL,

        -- Interruption Servicing
        PUSHF, POPF, RTI, LDISRA,

        -- Trap Servicing
        MFC, MFT, SYSCALL, LDTSRA

	);

	-- R8 processor instruction type. To be autogenerated by software
	--  Type 1 instructions are those which use regB as regBank(regTarget)
	--  Type 2 instructions are those which use regB as regBank(regSource2)
	--  Type 3 instructions are those which dont writeback to regBank
	type R8InstructionType_t is (Type1, Type2, Type3);

	-- Container for decoded instruction and its type
	type Instruction_t is record

		Instruction: R8Instruction_t;
		InstructionType: R8InstructionType_t;

	end record;

	-- State type for R8 processor state machine. To be autogenerated by software
	type State_t is (

		Sfetch, Sreg, Shalt, Sula, Swbk, Sld, Sst, Sjmp, Ssbrt, Spush, Srts, Spop, Sldsp,  -- Basic Instructions
		Smul, Sdiv, Smfh, Smfl,                                                            -- Multiplication and division
		Spushf, Spopf, Srti, Sitr, Sldisra,                                                -- Interruption servicing
		Sldtsra, Smfc, Smft, Ssyscall, Strap                                               -- Trap servicing
	);
    
	-- Decodes a given std_logic_vector to a R8 instruction and its type. To be autogenerated by software 
	function DecodeInstruction(InstructionValue: std_logic_vector(15 downto 0)) return Instruction_t;

	-- Defines processor registers as needed (e.g. defines regHIGH and regLOW only if multiplication and division should be supported). 
	--  To be auto generated by software.
	type ProcessorRegisters_t is record

		regPC    : std_logic_vector(15 downto 0);  -- Program Counter
		regIR    : std_logic_vector(15 downto 0);  -- Current Instruction (being executed)
		regSP    : std_logic_vector(15 downto 0);  -- Stack Pointer
        regALU   : std_logic_vector(15 downto 0);  -- ALU output register
        regA     : std_logic_vector(15 downto 0);  -- First reg bank output register
        regB     : std_logic_vector(15 downto 0);  -- Second reg bank output register
		regHIGH  : std_logic_vector(15 downto 0);  -- Higher order bits of multiplication result / division remainder
		regLOW   : std_logic_vector(15 downto 0);  -- Lower order bits of multiplication result / division quotient
        regISRA  : std_logic_vector(15 downto 0);  -- Address of Interruption Service Routine (ISR)
        regTSRA  : std_logic_vector(15 downto 0);  -- Address of Trap Service Routine (TSR)
        regCAUSE : std_logic_vector(15 downto 0);  -- Trap ID
        regITR   : std_logic_vector(15 downto 0);  -- Address of interruption/trap causing instruction

	end record;

	-- Declares processor registers
	signal ProcessorRegisters : ProcessorRegisters_t;
	alias regPC : std_logic_vector(15 downto 0) is ProcessorRegisters.regPC;
	alias regIR : std_logic_vector(15 downto 0) is ProcessorRegisters.regIR;
	alias regSP : std_logic_vector(15 downto 0) is ProcessorRegisters.regSP;
	

	-- All processor registers <= 0. To be autogenerated by software
	procedure ResetProcessorRegisters(ProcessorRegisters: inout ProcessorRegisters_t);

	-- Configuration values
	constant SupportsMultiplication: boolean := false;
	constant SupportsDivision: boolean := false;
	constant SupportsInterruptions: boolean := false;
	constant SupportsTraps: boolean := false;

	-- To be generated if multiplication is supported
	signal multiplicador: std_logic_vector(31 downto 0);

	-- To be generated if division is supported
	signal divisor: std_logic_vector(31 downto 0);



end package R8_PKG;


package body R8_PKG is


	-- Decodes a given std_logic_vector to a R8 instruction and its type. To be autogenerated by software 
	function DecodeInstruction(InstructionValue: std_logic_vector(15 downto 0)) return Instruction_t is

		-- Alias definitions for given instruction std_logic_vector
		alias OPCODE      : std_logic_vector(3 downto 0) is InstructionValue(15 downto 12);
		alias REGTARGET   : std_logic_vector(3 downto 0) is InstructionValue(11 downto 8);
		alias REGSOURCE1  : std_logic_vector(3 downto 0) is InstructionValue(7 downto 4);
		alias REGSOURCE2  : std_logic_vector(3 downto 0) is InstructionValue(3 downto 0);
		alias CONSTANTE   : std_logic_vector(7 downto 0) is InstructionValue(7 downto 0);
		alias JMPD_AUX    : std_logic_vector(1 downto 0) is InstructionValue(11 downto 10);
		alias JMPD_DESLOC : std_logic_vector(9 downto 0) is InstructionValue(9 downto 0);
		alias JSRD_DESLOC : std_logic_vector(11 downto 0) is InstructionValue(11 downto 0);

		-- Temp value for instruction and instruction type (to be returned)
		variable R8Instruction : Instruction_t;

	begin

		-- Decodes instruction
		if OPCODE = x"0" then R8instruction.Instruction := ADD; 
		elsif OPCODE = x"1" then R8instruction.Instruction := SUB;
		elsif OPCODE = x"2" then R8instruction.Instruction := AAND;
		elsif OPCODE = x"3" then R8instruction.Instruction := OOR;
		elsif OPCODE = x"4" then R8instruction.Instruction := XXOR;
		elsif OPCODE = x"5" then R8instruction.Instruction := ADDI;
		elsif OPCODE = x"6" then R8instruction.Instruction := SUBI;
		elsif OPCODE = x"7" then R8instruction.Instruction := LDL;
		elsif OPCODE = x"8" then R8instruction.Instruction := LDH;
		elsif OPCODE = x"9" then R8instruction.Instruction := LD;
		elsif OPCODE = x"A" then R8instruction.Instruction := ST;
		elsif OPCODE = x"B" and REGSOURCE2 = x"0" then R8instruction.Instruction := SL0;
		elsif OPCODE = x"B" and REGSOURCE2 = x"1" then R8instruction.Instruction := SL1;
		elsif OPCODE = x"B" and REGSOURCE2 = x"2" then R8instruction.Instruction := SR0;
		elsif OPCODE = x"B" and REGSOURCE2 = x"3" then R8instruction.Instruction := SR1;
		elsif OPCODE = x"B" and REGSOURCE2 = x"4" then R8instruction.Instruction := NNOT;
		elsif OPCODE = x"B" and REGSOURCE2 = x"5" then R8instruction.Instruction := NOP;
		elsif OPCODE = x"B" and REGSOURCE2 = x"6" then R8instruction.Instruction := HALT;
		elsif OPCODE = x"B" and REGSOURCE2 = x"7" then R8instruction.Instruction := LDSP;
		elsif OPCODE = x"B" and REGSOURCE2 = x"8" then R8instruction.Instruction := RTS;
		elsif OPCODE = x"B" and REGSOURCE2 = x"9" then R8instruction.Instruction := POP;
		elsif OPCODE = x"B" and REGSOURCE2 = x"A" then R8instruction.Instruction := PUSH;

		elsif OPCODE = x"B" and REGSOURCE2 = x"B" then R8instruction.Instruction := MUL;
		elsif OPCODE = x"B" and REGSOURCE2 = x"C" then R8instruction.Instruction := DIV;
		elsif OPCODE = x"B" and REGSOURCE2 = x"D" then R8instruction.Instruction := MFH;
		elsif OPCODE = x"B" and REGSOURCE2 = x"E" then R8instruction.Instruction := MFL;

		elsif OPCODE = x"B" and REGSOURCE2 = x"F" then R8instruction.Instruction := LDISRA;

		elsif OPCODE = x"C" and REGTARGET = x"0" and REGSOURCE2 = x"0" then R8instruction.Instruction := JMPR;
		elsif OPCODE = x"C" and REGTARGET = x"0" and REGSOURCE2 = x"1" then R8instruction.Instruction := JMPNR;
		elsif OPCODE = x"C" and REGTARGET = x"0" and REGSOURCE2 = x"2" then R8instruction.Instruction := JMPZR;
		elsif OPCODE = x"C" and REGTARGET = x"0" and REGSOURCE2 = x"3" then R8instruction.Instruction := JMPCR;
		elsif OPCODE = x"C" and REGTARGET = x"0" and REGSOURCE2 = x"4" then R8instruction.Instruction := JMPVR;

		elsif OPCODE = x"C" and REGTARGET = x"0" and REGSOURCE2 = x"5" then R8instruction.Instruction := JMP;
		elsif OPCODE = x"C" and REGTARGET = x"0" and REGSOURCE2 = x"6" then R8instruction.Instruction := JMPN;
		elsif OPCODE = x"C" and REGTARGET = x"0" and REGSOURCE2 = x"7" then R8instruction.Instruction := JMPZ;
		elsif OPCODE = x"C" and REGTARGET = x"0" and REGSOURCE2 = x"8" then R8instruction.Instruction := JMPC;
		elsif OPCODE = x"C" and REGTARGET = x"0" and REGSOURCE2 = x"9" then R8instruction.Instruction := JMPV;

		elsif OPCODE = x"D" and JMPD_AUX = "00" then R8instruction.Instruction := JMPD;
		elsif OPCODE = x"E" and JMPD_AUX = "00" then R8instruction.Instruction := JMPND;
		elsif OPCODE = x"E" and JMPD_AUX = "01" then R8instruction.Instruction := JMPZD;
		elsif OPCODE = x"E" and JMPD_AUX = "10" then R8instruction.Instruction := JMPCD;
		elsif OPCODE = x"E" and JMPD_AUX = "11" then R8instruction.Instruction := JMPVD;

		elsif OPCODE = x"C" and REGTARGET = x"0" and REGSOURCE2 = x"A" then R8instruction.Instruction := JSRR;
		elsif OPCODE = x"C" and REGTARGET = x"0" and REGSOURCE2 = x"B" then R8instruction.Instruction := JSR;
		elsif OPCODE = x"F" then R8instruction.Instruction := JSRD;

		elsif OPCODE = x"C" and REGTARGET = x"0" and REGSOURCE2 = x"C" then R8instruction.Instruction := PUSHF;
		elsif OPCODE = x"C" and REGTARGET = x"0" and REGSOURCE2 = x"D" then R8instruction.Instruction := POPF;
		elsif OPCODE = x"C" and REGTARGET = x"0" and REGSOURCE2 = x"E" then R8instruction.Instruction := RTI;

		elsif OPCODE = x"C" and REGTARGET = x"1" then R8instruction.Instruction := SYSCALL;
		elsif OPCODE = x"C" and REGTARGET = x"2" then R8instruction.Instruction := LDTSRA;
		elsif OPCODE = x"C" and REGTARGET = x"3" then R8instruction.Instruction := MFC;
		elsif OPCODE = x"C" and REGTARGET = x"4" then R8instruction.Instruction := MFT;

		else 

			R8instruction.Instruction := INVALID;
			report "INVALID instruction decoded" severity warning;

		end if;
		
		-- Decode instruction type
		if (R8instruction.Instruction = ADD or R8instruction.Instruction = SUB or R8instruction.Instruction = AAND or
           		R8instruction.Instruction = OOR  or R8instruction.Instruction = XXOR or R8instruction.Instruction = SL0 or
           		R8instruction.Instruction = SL1  or R8instruction.Instruction = SR0 or R8instruction.Instruction = SR1 or
           		R8instruction.Instruction = NOT_A) then

			R8Instruction.InstructionType = Type1;

        elsif (R8instruction.Instruction = ADDI or R8instruction.Instruction = SUBI or
              	R8instruction.Instruction = LDL  or R8instruction.Instruction = LDH) then

        	R8Instruction.InstructionType = Type2;

        else

        	R8Instruction.InstructionType = Type3;

        end if;

		return R8Instruction;
		
	end function DecodeInstruction;


	-- All processor registers <= 0. To be autogenerated by software
	procedure ResetProcessorRegisters(ProcessorRegisters : inout ProcessorRegisters_t) is begin

		-- Reset all processor registers (ProcessorRegisters_t is defined on package declaration)
		ProcessorRegisters.regPC    <= (others=>'0');
		ProcessorRegisters.regSP    <= (others=>'0');
        ProcessorRegisters.regALU   <= (others=>'0');
        ProcessorRegisters.regIR    <= (others=>'0');
        ProcessorRegisters.regA     <= (others=>'0');
        ProcessorRegisters.regB     <= (others=>'0');
		ProcessorRegisters.regFLAGS <= (others=>'0');
		ProcessorRegisters.regHIGH  <= (others=>'0');
		ProcessorRegisters.regLOW   <= (others=>'0');
        ProcessorRegisters.regISRA  <= (others=>'0');
        ProcessorRegisters.regTSRA  <= (others=>'0');
        ProcessorRegisters.regCAUSE <= (others=>'0');
        ProcessorRegisters.regITR   <= (others=>'0');
		
	end procedure ResetProcessorRegisters;


end package body R8_PKG;
